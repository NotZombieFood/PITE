import encoder_fec_pkg::*;

module encoder(
    input clk,
    input rst_n,
    input en,
    input message_data_t data_in,
    output encoded_message_data_t data_out
);


end module //encoder