import encoder_fec_pkg::*;

module decoder(
    input clk,
    input rst_n,
    input en,
    input demodulated_message_data_t data_in,
    output message_data_t data_out
);


end module //decoder